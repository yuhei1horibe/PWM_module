//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/05/2019 04:51:20 PM
// Design Name: 
// Module Name: PWM_UNIT_TEST
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifndef TRANS_GUARD
`define TRANS_GUARD

// Transaction generates patterns with constraints
// transaction is generated by generator.
class pwm_transaction;
    // Define transaction pattern
    rand bit [7:0] pwm_value;
    rand bit [7:0] pwm_range;

    constraint val_leq_range { pwm_value <= pwm_range; };
endclass

`endif
